module NOT_gate(input a, output out);
  assign out = ~a;
  //not n1(out,a);
endmodule
