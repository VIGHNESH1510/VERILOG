module OR_gate(input a,b,output out);
  assign out = a|b;
//   or o(out,a,b);
endmodule
