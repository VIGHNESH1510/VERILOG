module sathyan();

